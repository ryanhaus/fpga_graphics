typedef struct packed {
	integer x;
	integer y;
} point;

typedef struct packed {
	point a;
	point b;
	point c;
} triangle;
